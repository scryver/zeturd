tb_opcodes.vhd
